library verilog;
use verilog.vl_types.all;
entity tb_UART_TX is
end tb_UART_TX;
